library ieee;
use ieee.std_logic_1164.all;

package vga_640x480x1_frame_type is
        type vga_640x480x1_frame is array(0 to 640-1) of std_logic_vector(0 to 480-1);
end package;

package body vga_640x480x1_frame_type is
end package body vga_640x480x1_frame_type;
